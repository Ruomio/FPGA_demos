module clk (
    ports
);
    
endmodule